module demux_1X8();
	endmodule