module mux_8X1();
	endmodule