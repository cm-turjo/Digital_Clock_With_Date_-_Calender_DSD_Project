module breadboard();
	endmodule